module FOC();

endmodule