module iic_dri
#(
	parameter SLAVE_ADDR=7'b1010000,
	parameter CLK_FREQ  =26'd50_000_000,
	parameter IIC_FREQ  =28'd250_000
)(
	input clk,
	input rst_n,
	//iic interface
	input 				iic_exec,
	input 				bit_ctrl,
	input 				iic_rh_wl,
	input[15:0] 		iic_addr,
	input[7:0]			iic_data_w,
	output reg[7:0]	iic_data_r,
	output reg			iic_done,
	output reg			scl,
	inout					sda,
	output reg			dri_clk
);
//parameters
localparam	IDLE		='b0000_0001;
localparam	SLADDR	='b0000_0001;
localparam	ADDRL		='b0000_0001;
localparam	ADDRH		='b0000_0001;
localparam	DATA_WR	='b0000_0001;
localparam	ADDR_RD	='b0000_0001;
localparam	DATA_RD	='b0000_0001;
localparam	STOP		='b0000_0001;
//registers
reg 			sda_dir;
reg 			sda_out;
reg 			wr_flag;
reg 			st_done;
reg[6:0] 	cnt;
reg[7:0] 	cur_state;
reg[7:0] 	next_state;
reg[15:0]	addr_t;
reg[7:0] 	data_r;
reg[7:0] 	data_wr_t;
reg[9:0] 	clk_cnt;
//wires
wire 			sda_in;
wire[8:0]	clk_divide;

assign sda			=sda_dir ? sda_out : 1'bz;
assign sda_in		=sda;
assign clk_divide	=(CLK_FREQ/IIC_FREQ)>>2'd3;
always @(posedge clk or negedge rst_n)begin
	if(!rst_n) begin
        dri_clk <=  1'b1;
        clk_cnt <= 10'd0;
    end
    else if(clk_cnt == clk_divide - 1'd1) begin
        clk_cnt <= 10'd0;
        dri_clk <= ~dri_clk;	//此为1MHz，后面操作时还会再4分频
    end
    else
        clk_cnt <= clk_cnt + 1'b1;
end
//(三段式状态机)同步时序描述状态转移
always @(posedge dri_clk or negedge rst_n) begin
    if(!rst_n)
        cur_state <= IDLE;
    else
        cur_state <= next_state;
end

//组合逻辑判断状态转移条件
always @( * ) begin
//    next_state = st_idle;
    case(cur_state)
        IDLE: begin                            // 空闲状态
           if(iic_exec) begin	//如果有触发信号
               next_state = SLADDR;
           end
           else
               next_state = IDLE;
        end
        SLADDR: begin
            if(st_done) begin
                if(bit_ctrl)                      // 判断是16位还是8位字地址
                   next_state = ADDRL;
                else
                   next_state = ADDRH ;
            end
            else
                next_state = SLADDR;
        end
        ADDRL: begin                          // 写16位字地址
            if(st_done) begin
                next_state = ADDRH;
            end
            else begin
                next_state = ADDRL;
            end
        end
        ADDRH: begin                           // 8位字地址
            if(st_done) begin
                if(!wr_flag)                 // 读写判断
                    next_state = DATA_WR;
                else
                    next_state = ADDR_RD;
            end
            else begin
                next_state = ADDRH;
            end
        end
        DATA_WR: begin                        // 写数据(8 bit)
            if(st_done)
                next_state = STOP;
            else
                next_state = DATA_WR;
        end
        ADDR_RD: begin                         // 写地址以进行读数据
            if(st_done) begin
                next_state = DATA_RD;
            end
            else begin
                next_state = ADDR_RD;
            end
        end
        DATA_RD: begin                        // 读取数据(8 bit)
            if(st_done)
                next_state = STOP;
            else
                next_state = DATA_RD;
        end
        STOP: begin                           // 结束iic操作
            if(st_done)
                next_state = IDLE;
            else
                next_state = STOP ;
        end
        default: next_state= IDLE;
    endcase
end
//时序电路描述状态输出
always @(posedge dri_clk or negedge rst_n) begin		//1MHz的时钟频率触发
    //复位初始化
    if(!rst_n) begin
        scl        <= 1'b1;
        sda_out    <= 1'b1;
        sda_dir    <= 1'b1;
        iic_done   <= 1'b0;
        cnt        <= 1'b0;
        st_done    <= 1'b0;
        data_r     <= 1'b0;
        iic_data_r <= 1'b0;
        wr_flag    <= 1'b0;
        addr_t     <= 1'b0;
        data_wr_t  <= 1'b0;
    end
    else begin
        st_done <= 1'b0 ;
        cnt     <= cnt +1'b1 ;	//计数自加，用于时序步骤递增
        case(cur_state)	//判断当前状态
            IDLE: begin                             // 空闲状态
                scl     <= 1'b1;	// IIC协议规定，时钟线和数据线均为高时，代表空闲
                sda_out <= 1'b1;
                sda_dir <= 1'b1;	// sda为输出模式，
                iic_done<= 1'b0;
                cnt     <= 7'b0;
                if(iic_exec) begin
                    wr_flag   <= iic_rh_wl ;			//读写信号
                    addr_t    <= iic_addr  ;			//iic器件内地址
                    data_wr_t <= iic_data_w;			//需要写入的数据
                end
            end
            SLADDR: begin                            // 写器件地址和“写”信号
                case(cnt)
                    7'd1 : sda_out <= 1'b0;             // 开始iic，参考IIC协议时序图
                    7'd3 : scl <= 1'b0;					
                    7'd4 : sda_out <= SLAVE_ADDR[6];    // 传送器件地址
                    7'd5 : scl <= 1'b1;  
                    7'd7 : scl <= 1'b0;//此处scl的高低电平变化为每4个时钟一个周期，即250KHz，因此跳过6
                    7'd8 : sda_out <= SLAVE_ADDR[5];
                    7'd9 : scl <= 1'b1;
                    7'd11: scl <= 1'b0;
                    7'd12: sda_out <= SLAVE_ADDR[4];
                    7'd13: scl <= 1'b1;
                    7'd15: scl <= 1'b0;
                    7'd16: sda_out <= SLAVE_ADDR[3];
                    7'd17: scl <= 1'b1;
                    7'd19: scl <= 1'b0;
                    7'd20: sda_out <= SLAVE_ADDR[2];
                    7'd21: scl <= 1'b1;
                    7'd23: scl <= 1'b0;
                    7'd24: sda_out <= SLAVE_ADDR[1];
                    7'd25: scl <= 1'b1;
                    7'd27: scl <= 1'b0;
                    7'd28: sda_out <= SLAVE_ADDR[0];
                    7'd29: scl <= 1'b1;
                    7'd31: scl <= 1'b0;
                    7'd32: sda_out <= 1'b0;              // 0:写
                    7'd33: scl <= 1'b1;
                    7'd35: scl <= 1'b0;
                    7'd36: begin
                        sda_dir <= 1'b0;                 // sda变为高阻态
                        sda_out <= 1'b1;				 // 拉高sda，等待从机应答
                    end
                    7'd37: scl     <= 1'b1;
                    7'd38: st_done <= 1'b1;				 // 一个状态结束信号
                    7'd39: begin
                        scl <= 1'b0;
                        cnt <= 1'b0;
                    end
                    default :  ;
                endcase
            end
            ADDRL: begin
                case(cnt)
                    7'd0 : begin
                        sda_dir <= 1'b1 ;
                        sda_out <= addr_t[15];           // 传送内地址的高8位
                    end
                    7'd1 : scl <= 1'b1;
                    7'd3 : scl <= 1'b0;
                    7'd4 : sda_out <= addr_t[14];
                    7'd5 : scl <= 1'b1;
                    7'd7 : scl <= 1'b0;
                    7'd8 : sda_out <= addr_t[13];
                    7'd9 : scl <= 1'b1;
                    7'd11: scl <= 1'b0;
                    7'd12: sda_out <= addr_t[12];
                    7'd13: scl <= 1'b1;
                    7'd15: scl <= 1'b0;
                    7'd16: sda_out <= addr_t[11];
                    7'd17: scl <= 1'b1;
                    7'd19: scl <= 1'b0;
                    7'd20: sda_out <= addr_t[10];
                    7'd21: scl <= 1'b1;
                    7'd23: scl <= 1'b0;
                    7'd24: sda_out <= addr_t[9];
                    7'd25: scl <= 1'b1;
                    7'd27: scl <= 1'b0;
                    7'd28: sda_out <= addr_t[8];
                    7'd29: scl <= 1'b1;
                    7'd31: scl <= 1'b0;
                    7'd32: begin
                        sda_dir <= 1'b0;                 // 从机应答
                        sda_out <= 1'b1;
                    end
                    7'd33: scl     <= 1'b1;
                    7'd34: st_done <= 1'b1;
                    7'd35: begin
                        scl <= 1'b0;
                        cnt <= 1'b0;
                    end
                    default :  ;
                endcase
            end
            ADDRH: begin
                case(cnt)
                    7'd0: begin
                       sda_dir <= 1'b1 ;
                       sda_out <= addr_t[7];            // 16位时传输内地址的低8位，8位时传送8位地址
                    end
                    7'd1 : scl <= 1'b1;
                    7'd3 : scl <= 1'b0;
                    7'd4 : sda_out <= addr_t[6];
                    7'd5 : scl <= 1'b1;
                    7'd7 : scl <= 1'b0;
                    7'd8 : sda_out <= addr_t[5];
                    7'd9 : scl <= 1'b1;
                    7'd11: scl <= 1'b0;
                    7'd12: sda_out <= addr_t[4];
                    7'd13: scl <= 1'b1;
                    7'd15: scl <= 1'b0;
                    7'd16: sda_out <= addr_t[3];
                    7'd17: scl <= 1'b1;
                    7'd19: scl <= 1'b0;
                    7'd20: sda_out <= addr_t[2];
                    7'd21: scl <= 1'b1;
                    7'd23: scl <= 1'b0;
                    7'd24: sda_out <= addr_t[1];
                    7'd25: scl <= 1'b1;
                    7'd27: scl <= 1'b0;
                    7'd28: sda_out <= addr_t[0];
                    7'd29: scl <= 1'b1;
                    7'd31: scl <= 1'b0;
                    7'd32: begin
                        sda_dir <= 1'b0;                // 从机应答
                        sda_out <= 1'b1;
                    end
                    7'd33: scl     <= 1'b1;
                    7'd34: st_done <= 1'b1;
                    7'd35: begin
                        scl <= 1'b0;
                        cnt <= 1'b0;
                    end
                    default :  ;
                endcase
            end
            DATA_WR: begin                          // 写数据(8 bit)
                case(cnt)
                    7'd0: begin
                        sda_out <= data_wr_t[7];        // iic写8位数据
                        sda_dir <= 1'b1;
                    end
                    7'd1 : scl <= 1'b1;
                    7'd3 : scl <= 1'b0;
                    7'd4 : sda_out <= data_wr_t[6];
                    7'd5 : scl <= 1'b1;
                    7'd7 : scl <= 1'b0;
                    7'd8 : sda_out <= data_wr_t[5];
                    7'd9 : scl <= 1'b1;
                    7'd11: scl <= 1'b0;
                    7'd12: sda_out <= data_wr_t[4];
                    7'd13: scl <= 1'b1;
                    7'd15: scl <= 1'b0;
                    7'd16: sda_out <= data_wr_t[3];
                    7'd17: scl <= 1'b1;
                    7'd19: scl <= 1'b0;
                    7'd20: sda_out <= data_wr_t[2];
                    7'd21: scl <= 1'b1;
                    7'd23: scl <= 1'b0;
                    7'd24: sda_out <= data_wr_t[1];
                    7'd25: scl <= 1'b1;
                    7'd27: scl <= 1'b0;
                    7'd28: sda_out <= data_wr_t[0];
                    7'd29: scl <= 1'b1;
                    7'd31: scl <= 1'b0;
                    7'd32: begin
                        sda_dir <= 1'b0;                // 从机应答
                        sda_out <= 1'b1;
                    end
                    7'd33: scl <= 1'b1;
                    7'd34: st_done <= 1'b1;
                    7'd35: begin
                        scl  <= 1'b0;
                        cnt  <= 1'b0;
                    end
                    default  :  ;
                endcase
            end
            ADDR_RD: begin                           // 写器件地址和“读”信号以进行读数据
                case(cnt)
                    7'd0 : begin
                        sda_dir <= 1'b1;
                        sda_out <= 1'b1;
                    end
                    7'd1 : scl <= 1'b1;
                    7'd2 : sda_out <= 1'b0;             // 重新开始
                    7'd3 : scl <= 1'b0;
                    7'd4 : sda_out <= SLAVE_ADDR[6];    // 传送器件地址
                    7'd5 : scl <= 1'b1;
                    7'd7 : scl <= 1'b0;
                    7'd8 : sda_out <= SLAVE_ADDR[5];
                    7'd9 : scl <= 1'b1;
                    7'd11: scl <= 1'b0;
                    7'd12: sda_out <= SLAVE_ADDR[4];
                    7'd13: scl <= 1'b1;
                    7'd15: scl <= 1'b0;
                    7'd16: sda_out <= SLAVE_ADDR[3];
                    7'd17: scl <= 1'b1;
                    7'd19: scl <= 1'b0;
                    7'd20: sda_out <= SLAVE_ADDR[2];
                    7'd21: scl <= 1'b1;
                    7'd23: scl <= 1'b0;
                    7'd24: sda_out <= SLAVE_ADDR[1];
                    7'd25: scl <= 1'b1;
                    7'd27: scl <= 1'b0;
                    7'd28: sda_out <= SLAVE_ADDR[0];
                    7'd29: scl <= 1'b1;
                    7'd31: scl <= 1'b0;
                    7'd32: sda_out <= 1'b1;             // 1:读
                    7'd33: scl <= 1'b1;
                    7'd35: scl <= 1'b0;
                    7'd36: begin
                        sda_dir <= 1'b0;                // 从机应答
                        sda_out <= 1'b1;
                    end
                    7'd37: scl     <= 1'b1;
                    7'd38: st_done <= 1'b1;
                    7'd39: begin
                        scl <= 1'b0;
                        cnt <= 1'b0;
                    end
                    default : ;
                endcase
            end
            DATA_RD: begin                          // 读取数据(8 bit)
                case(cnt)
                    7'd0: sda_dir <= 1'b0;			   // sda高阻态，等待读数据
                    7'd1: begin
                        data_r[7] <= sda_in;
                        scl       <= 1'b1;
                    end
                    7'd3: scl  <= 1'b0;
                    7'd5: begin
                        data_r[6] <= sda_in ;
                        scl       <= 1'b1   ;
                    end
                    7'd7: scl  <= 1'b0;
                    7'd9: begin
                        data_r[5] <= sda_in;
                        scl       <= 1'b1  ;
                    end
                    7'd11: scl  <= 1'b0;
                    7'd13: begin
                        data_r[4] <= sda_in;
                        scl       <= 1'b1  ;
                    end
                    7'd15: scl  <= 1'b0;
                    7'd17: begin
                        data_r[3] <= sda_in;
                        scl       <= 1'b1  ;
                    end
                    7'd19: scl  <= 1'b0;
                    7'd21: begin
                        data_r[2] <= sda_in;
                        scl       <= 1'b1  ;
                    end
                    7'd23: scl  <= 1'b0;
                    7'd25: begin
                        data_r[1] <= sda_in;
                        scl       <= 1'b1  ;
                    end
                    7'd27: scl  <= 1'b0;
                    7'd29: begin
                        data_r[0] <= sda_in;
                        scl       <= 1'b1  ;
                    end
                    7'd31: scl  <= 1'b0;
                    7'd32: begin
                        sda_dir <= 1'b1;              // sda输出，将由主机给出是否应答
                        sda_out <= 1'b1;			  // 主机将sda拉高，表示非应答，结束本次读取
                    end
                    7'd33: scl     <= 1'b1;
                    7'd34: st_done <= 1'b1;
                    7'd35: begin
                        scl <= 1'b0;
                        cnt <= 1'b0;
                        iic_data_r <= data_r;
                    end
                    default  :  ;
                endcase
            end
            STOP: begin                            // 结束iic操作
                case(cnt)
                    7'd0: begin
                        sda_dir <= 1'b1;              // 结束iic
                        sda_out <= 1'b0;
                    end
                    7'd1 : scl     <= 1'b1;
                    7'd3 : sda_out <= 1'b1;
                    7'd15: st_done <= 1'b1;
                    7'd16: begin
                        cnt      <= 1'b0;
                        iic_done <= 1'b1;             // 向上层模块传递iic结束信号
                    end
                	default  : ;
                endcase
            end
        endcase
    end
end

endmodule
